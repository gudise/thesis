`define LOW 2'b00
`define RISING 2'b01
`define FALLING 2'b10
`define HIGH 2'b11

`define IDLE        1
`define RST         2
`define RST_SYNC    3
`define CALC        4
`define CALC_SYNC   5
`define SCAN        6
`define SCAN_SYNC   7
`define PRINT       8
`define PRINT_SYNC  9

`define cmd_idle        0
`define cmd_reset       1
`define cmd_calc        2
`define cmd_scan        3
`define cmd_print       4
`define cmd_end	        5

`define cmd_idle_sync	 6
`define cmd_reset_sync	 7
`define cmd_calc_sync	 8
`define cmd_scan_sync    9
`define cmd_print_sync   10
