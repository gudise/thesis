/*
 Este módulo implementa una interfaz para conectar el sistema de procesamiento (PS/MicroBlaze) con la lógica
 programable de la FPGA (PL). La forma de comunicarse con PS es a través de una máquina de estados (FSM) que
 es controlada por PS mediante un canal 'ctrl', de acuerdo con un cierto protocolo. La comunicación con PL 
 se hace a través de un protocolo 'handshake', de modo que cuando la interfaz dispone de un dato disponible
 sube una señal 'sync'->1; una vez los cálculos en PL han terminado, la interfaz espera recibir 'ack'->1. Por
 último, para reiniciar el ciclo de lectura, la interfaz bajará 'sync'->0, y cuando reciba 'ack'->0 proseguirá
 la comunicación con PS. 
*/

`include "interfaz_pspl_define.vh"


`define LOW		2'b00
`define RISING	2'b01
`define FALLING	2'b10
`define HIGH	2'b11

`define IDLE		1
`define CALC		2
`define CALC_SYNC	3
`define SCAN		4
`define SCAN_SYNC	5
`define PRINT		6
`define PRINT_SYNC	7

`define cmd_idle		0
`define cmd_calc		1
`define cmd_scan		2
`define cmd_print		3
`define cmd_end			4
`define cmd_idle_sync	5
`define cmd_calc_sync	6
`define cmd_scan_sync	7
`define cmd_print_sync	8

module INTERFAZ_PSPL #(
	parameter	DATA_WIDTH=32,
	parameter	BUFFER_IN_WIDTH=16,
	parameter	BUFFER_OUT_WIDTH=16
	) (
	input							clock,
	input[7:0]						ctrl_in,	// instrucción de PS.
	output reg[7:0]					ctrl_out,	// instrucción a PS.
	input[DATA_WIDTH-1:0]			data_in,	// dato de PS.
	output reg[DATA_WIDTH-1:0]		data_out,	// dato a PS.
	output reg						sync=0,		//
	input							ack,		// intefaz 'handshake' con PL.
	output reg[BUFFER_IN_WIDTH-1:0]	buffer_in,	// 'buffer' enviado por PS.
	input[BUFFER_OUT_WIDTH-1:0]		buffer_out	// 'buffer' devuelto a PS.
	);

	reg[3:0] state=`IDLE;
	reg[1:0] busy_frontend=`LOW;
	reg[1:0] busy_backend=`LOW;
	reg[7:0] ctrl_in_reg;
	reg[DATA_WIDTH-1:0] data_in_reg;
	reg[7:0] contador_std;
	
	//registro de input
	always @(posedge clock) begin
		ctrl_in_reg <= ctrl_in;
		data_in_reg <= data_in;
	end
	 
	//definicion de estados
	always @(posedge clock) begin
		busy_frontend[1] <= busy_frontend[0];
		case (state)
			`IDLE: begin
				//condicion de estabilidad de 'IDLE'
				if(!sync && !ack) busy_frontend[0] <= 1;
				else busy_frontend[0] <= 0;
				
				sync <= 0;
			end
			
			`CALC: begin
				//condicion de estabilidad de 'CALC'
				if(ack) busy_frontend[0] <= 1;
				else busy_frontend[0] <= 0;
				
				sync <= 1;
			end
		endcase
	end

	//bucle dinamico estandar
	always @(posedge clock) begin
		busy_backend[1] <= busy_backend[0];  
		case(state)

			`IDLE: begin
				ctrl_out <= `cmd_idle_sync;
				
				contador_std <= 0;
				
				case(ctrl_in_reg)
					`cmd_calc: begin
						state <= `CALC;
						busy_backend[0] <= 0;
					end
					`cmd_scan: begin
						state <= `SCAN;
						busy_backend[0] <= 0;
					end
					`cmd_print: begin
						state <= `PRINT;
						busy_backend[0] <= 0;
					end
					default: begin
						state <= `IDLE;
						busy_backend[0] <= 1;
					end
				endcase
			end
			
			`CALC: begin
				if(busy_frontend==`HIGH && busy_backend==`HIGH) begin
					state <= `CALC_SYNC;
					busy_backend[0] <= 0;
				end
				else begin
					state <= `CALC;
					busy_backend[0] <= 1;
				end				
			end
			
			`CALC_SYNC: begin
				ctrl_out <= `cmd_calc_sync;
				
				if(ctrl_in_reg==`cmd_idle) begin
					state <= `IDLE;
					busy_backend[0] <= 0;
				end
				else begin
					state <= `CALC_SYNC;
					busy_backend[0] <= 1;
				end
			end
			
			`SCAN: begin
				ctrl_out <= `cmd_scan;
				
				if(ctrl_in_reg==`cmd_scan_sync) begin
					`ifdef DW_GT_BIW
						buffer_in <= data_in;
					
					`elsif BIW_ALIGNED_DW
						buffer_in[DATA_WIDTH*(contador_std+1)-1 -: DATA_WIDTH] <= data_in;
						
					`elsif BIW_MISALIGNED_DW
						if(contador_std<BUFFER_IN_WIDTH/DATA_WIDTH)
							buffer_in[DATA_WIDTH*(contador_std+1)-1 -: DATA_WIDTH] <= data_in;
						else if(contador_std==BUFFER_IN_WIDTH/DATA_WIDTH)
							buffer_in[BUFFER_IN_WIDTH-1 : BUFFER_IN_WIDTH-BUFFER_IN_WIDTH%DATA_WIDTH] <= data_in;
							
					`else
						buffer_in <= data_in;
						
					`endif
					
					state <= `SCAN_SYNC;
					busy_backend[0] <= 0;
				end
				else begin
					state <= `SCAN;
					busy_backend[0] <= 1;
				end
			end
			
			`SCAN_SYNC: begin
				ctrl_out <= `cmd_scan_sync;
				
				if(ctrl_in_reg==`cmd_idle) begin
					state <= `IDLE;
					busy_backend[0] <= 0;
				end
				else if(ctrl_in_reg==`cmd_scan) begin
					state <= `SCAN;
					contador_std <= contador_std + 1;
					busy_backend[0] <= 0;
				end
				else begin
					state <= `SCAN_SYNC;
					busy_backend[0] <= 1;
				end
			end
			
			`PRINT: begin
				ctrl_out <= `cmd_print;
								
				`ifdef DW_GT_BOW
					data_out <= buffer_out;
					
				`elsif BOW_ALIGNED_DW
					data_out <= buffer_out[DATA_WIDTH*(contador_std+1)-1 -: DATA_WIDTH];
				
				`elsif BOW_MISALIGNED_DW
					if(contador_std<BUFFER_OUT_WIDTH/DATA_WIDTH)
						data_out <= buffer_out[DATA_WIDTH*(contador_std+1)-1 -: DATA_WIDTH];
					else if(contador_std==BUFFER_OUT_WIDTH/DATA_WIDTH)
						data_out <= buffer_out[BUFFER_OUT_WIDTH-1 : BUFFER_OUT_WIDTH-BUFFER_OUT_WIDTH%DATA_WIDTH];
				
				`else
					data_out <= buffer_out;
				
				`endif
				
				if(ctrl_in_reg==`cmd_print_sync) begin
					state <= `PRINT_SYNC;
					busy_backend[0] <= 0;
				end
				else begin
					state <= `PRINT;
					busy_backend[0] <= 1;
				end
			end
			
			`PRINT_SYNC: begin
				ctrl_out <= `cmd_print_sync;
								
				if(ctrl_in_reg==`cmd_idle) begin
					state <= `IDLE;
					busy_backend[0] <= 0;
				end
				else if(ctrl_in_reg==`cmd_print) begin
					state <= `PRINT;
					contador_std <= contador_std + 1;
					busy_backend[0] <= 0;
				end
				else begin
					state <= `PRINT_SYNC;
					busy_backend[0] <= 1;
				end
			end
		endcase
	end

endmodule
